interface dff_Interface();
  logic [7:0] din;
  logic rst;
  logic clk;
  logic [7:0] dout;
endinterface